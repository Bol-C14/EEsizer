* RC lowpass example (no .control)
V1 in 0 AC 1
R1 in out 10k
C1 out 0 1u
Rleak out 0 1G
.end
