* RC lowpass example (no .control)
V1 in 0 AC 1
R1 in out 1k
C1 out 0 1u
.end
